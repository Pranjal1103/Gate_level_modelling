module not_g(y,a);
  input a;
  output y;
  not n1(y,a);
endmodule
