module nand_g(y,a,b);
  input a,b;
  output y;
  nand n1(y,a,b);
endmodule
