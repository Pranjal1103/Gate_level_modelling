module or_g(y,a,b);
  input a,b;
  output y;
  or n1(y,a,b);
endmodule
