module xor_g(y,a,b);
  input a,b;
  output y;
  xor n1(y,a,b);
endmodule
