module nor_g(y,a,b);
  input a,b;
  output y;
  nor n1(y,a,b);
endmodule
