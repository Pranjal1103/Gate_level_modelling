module and_g(y,a,b);
  input a,b;
  output y;
  and n1(y,a,b);
endmodule
